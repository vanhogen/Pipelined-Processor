module or2(inA, inB, Out);
    input inA;
    input inB;
    output Out;
    assign Out = inA | inB;
endmodule
